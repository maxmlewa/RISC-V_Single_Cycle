`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: imm_gen
// Project Name: Single Cycle Processor
// Target Devices: XXXX
// Description: Immediate Generator for RV32I instructions
//              Extracts and sign-extends immediate fields from 32 bit instruction
//              Operation based on the instruction format: I, S, B, U, J
// 
// Dependencies: None, pure standalone module
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module imm_gen(

    );
endmodule
