`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////

// Module Name: instr_memory
// Project Name: Single Cycle Processor
// Target Devices: XXXX
// Description: Instruction Memory for the RV32I Single Cycle Processor
//              Single read port that performs a combinational read 
//              Not clocked, because the memory has no write port
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module instr_memory(

    );
endmodule
