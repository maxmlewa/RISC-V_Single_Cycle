`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: regfile
// Project Name: Single Cycle Processor
// Target Devices: XXXX
// Description: Register File for RV321
//              2 read ports and 1 write port
//              Synchronous write and asynchronous reads
// 
// Dependencies: No defined modules instantiated
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module regfile(

    );
endmodule
