`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: testbench_imm_gen
// Project Name: 
// Target Devices:
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_imm_gen(

    );
endmodule
