`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Module Name: testbench_alu
// Project Name: Single Cycle Processor
// Target Devices: XXXX
// Description: Unit testbench for the alu module
// 
// Dependencies: alu.v: alu module instantiated as the DUT
// Functionality tested: ADD, SUB, SLT, SLTU, AND, OR, XOR, SLL, SRL, SRA
//                       Proper ALU control signal decoding from instruction fields
//                       Zero output flag for branch comparisons
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module testbench_alu( );
    
    // 
endmodule
