`timescale 1ns / 1ps
////////////////////////////////////////////////////////////////////////////////// 
// Module Name: control_unit
// Project Name: Single Cycle Processor
// Target Devices: XXXX
// Description: Main control logic for RV32I
//              Decodes the opcode (and funct3 for the memory access width)
//              Generates the control signals for the datapath component
// 
// Dependencies: None, pure standalone
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module control_unit(

    );
endmodule
